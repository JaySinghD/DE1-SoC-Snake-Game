
//General item spawn that will work for apples or powerups
module itemSpawn(input CLOCK_50, input [3:0] snakePositionX, input [3:0] snakePositionY, output reg [3:0] spawnPositionX, output reg [3:0] spawnPositionY,output reg [7:0] snakeLength, output reg [1:0] gameClockSelect, output reg [2:0] itemColour);
   
   //takes in itemEaten, which signifies that if the item needs to be replaced
   
   //outputs newItemEaten, which signifies that the item.
   
  
   // input itemEaten;

    reg [7:0] xySelector; //256 different values, from 0 to 255,,,,, must stop after 224

    reg [3:0] grid_x [0:224];
    reg [3:0] grid_y [0:224];

    //fills in the appropriate square
    //fillGridSq square(spawnPositionX, spawnPositionY, clr, 1'b1, CLOCK_50);

    initial begin
        //statements to execute once
        xySelector = 8'd0;
        snakeLength = 1;

        //Defining all positions -> Generated by ChatGPT
        grid_x[0] = 4'd2; grid_y[0] = 4'd8;
        grid_x[1] = 4'd14; grid_y[1] = 4'd3;
        grid_x[2] = 4'd10; grid_y[2] = 4'd11;
        grid_x[3] = 4'd8; grid_y[3] = 4'd14;
        grid_x[4] = 4'd9; grid_y[4] = 4'd5;
        grid_x[5] = 4'd4; grid_y[5] = 4'd14;
        grid_x[6] = 4'd4; grid_y[6] = 4'd0;
        grid_x[7] = 4'd11; grid_y[7] = 4'd6;
        grid_x[8] = 4'd10; grid_y[8] = 4'd2;
        grid_x[9] = 4'd0; grid_y[9] = 4'd3;
        grid_x[10] = 4'd8; grid_y[10] = 4'd1;
        grid_x[11] = 4'd13; grid_y[11] = 4'd6;
        grid_x[12] = 4'd12; grid_y[12] = 4'd3;
        grid_x[13] = 4'd14; grid_y[13] = 4'd1;
        grid_x[14] = 4'd13; grid_y[14] = 4'd13;
        grid_x[15] = 4'd11; grid_y[15] = 4'd1;
        grid_x[16] = 4'd6; grid_y[16] = 4'd7;
        grid_x[17] = 4'd1; grid_y[17] = 4'd1;
        grid_x[18] = 4'd12; grid_y[18] = 4'd4;
        grid_x[19] = 4'd9; grid_y[19] = 4'd12;
        grid_x[20] = 4'd11; grid_y[20] = 4'd11;
        grid_x[21] = 4'd11; grid_y[21] = 4'd12;
        grid_x[22] = 4'd2; grid_y[22] = 4'd10;
        grid_x[23] = 4'd6; grid_y[23] = 4'd14;
        grid_x[24] = 4'd14; grid_y[24] = 4'd11;
        grid_x[25] = 4'd11; grid_y[25] = 4'd3;
        grid_x[26] = 4'd3; grid_y[26] = 4'd12;
        grid_x[27] = 4'd9; grid_y[27] = 4'd4;
        grid_x[28] = 4'd11; grid_y[28] = 4'd0;
        grid_x[29] = 4'd9; grid_y[29] = 4'd7;
        grid_x[30] = 4'd5; grid_y[30] = 4'd11;
        grid_x[31] = 4'd6; grid_y[31] = 4'd9;
        grid_x[32] = 4'd4; grid_y[32] = 4'd13;
        grid_x[33] = 4'd9; grid_y[33] = 4'd14;
        grid_x[34] = 4'd2; grid_y[34] = 4'd4;
        grid_x[35] = 4'd6; grid_y[35] = 4'd8;
        grid_x[36] = 4'd7; grid_y[36] = 4'd7;
        grid_x[37] = 4'd2; grid_y[37] = 4'd11;
        grid_x[38] = 4'd8; grid_y[38] = 4'd13;
        grid_x[39] = 4'd3; grid_y[39] = 4'd13;
        grid_x[40] = 4'd13; grid_y[40] = 4'd7;
        grid_x[41] = 4'd4; grid_y[41] = 4'd6;
        grid_x[42] = 4'd4; grid_y[42] = 4'd8;
        grid_x[43] = 4'd2; grid_y[43] = 4'd1;
        grid_x[44] = 4'd2; grid_y[44] = 4'd6;
        grid_x[45] = 4'd8; grid_y[45] = 4'd0;
        grid_x[46] = 4'd12; grid_y[46] = 4'd7;
        grid_x[47] = 4'd12; grid_y[47] = 4'd11;
        grid_x[48] = 4'd11; grid_y[48] = 4'd7;
        grid_x[49] = 4'd9; grid_y[49] = 4'd11;
        grid_x[50] = 4'd7; grid_y[50] = 4'd10;
        grid_x[51] = 4'd7; grid_y[51] = 4'd5;
        grid_x[52] = 4'd8; grid_y[52] = 4'd6;
        grid_x[53] = 4'd9; grid_y[53] = 4'd0;
        grid_x[54] = 4'd14; grid_y[54] = 4'd10;
        grid_x[55] = 4'd7; grid_y[55] = 4'd8;
        grid_x[56] = 4'd11; grid_y[56] = 4'd8;
        grid_x[57] = 4'd11; grid_y[57] = 4'd2;
        grid_x[58] = 4'd13; grid_y[58] = 4'd8;
        grid_x[59] = 4'd14; grid_y[59] = 4'd2;
        grid_x[60] = 4'd1; grid_y[60] = 4'd7;
        grid_x[61] = 4'd8; grid_y[61] = 4'd5;
        grid_x[62] = 4'd3; grid_y[62] = 4'd2;
        grid_x[63] = 4'd6; grid_y[63] = 4'd5;
        grid_x[64] = 4'd8; grid_y[64] = 4'd9;
        grid_x[65] = 4'd5; grid_y[65] = 4'd14;
        grid_x[66] = 4'd9; grid_y[66] = 4'd9;
        grid_x[67] = 4'd3; grid_y[67] = 4'd5;
        grid_x[68] = 4'd12; grid_y[68] = 4'd10;
        grid_x[69] = 4'd7; grid_y[69] = 4'd13;
        grid_x[70] = 4'd14; grid_y[70] = 4'd12;
        grid_x[71] = 4'd3; grid_y[71] = 4'd11;
        grid_x[72] = 4'd8; grid_y[72] = 4'd10;
        grid_x[73] = 4'd5; grid_y[73] = 4'd9;
        grid_x[74] = 4'd10; grid_y[74] = 4'd4;
        grid_x[75] = 4'd4; grid_y[75] = 4'd1;
        grid_x[76] = 4'd12; grid_y[76] = 4'd8;
        grid_x[77] = 4'd1; grid_y[77] = 4'd13;
        grid_x[78] = 4'd4; grid_y[78] = 4'd9;
        grid_x[79] = 4'd13; grid_y[79] = 4'd2;
        grid_x[80] = 4'd14; grid_y[80] = 4'd4;
        grid_x[81] = 4'd11; grid_y[81] = 4'd10;
        grid_x[82] = 4'd8; grid_y[82] = 4'd8;
        grid_x[83] = 4'd0; grid_y[83] = 4'd5;
        grid_x[84] = 4'd7; grid_y[84] = 4'd4;
        grid_x[85] = 4'd13; grid_y[85] = 4'd5;
        grid_x[86] = 4'd3; grid_y[86] = 4'd3;
        grid_x[87] = 4'd5; grid_y[87] = 4'd6;
        grid_x[88] = 4'd13; grid_y[88] = 4'd4;
        grid_x[89] = 4'd8; grid_y[89] = 4'd3;
        grid_x[90] = 4'd13; grid_y[90] = 4'd10;
        grid_x[91] = 4'd2; grid_y[91] = 4'd5;
        grid_x[92] = 4'd0; grid_y[92] = 4'd12;
        grid_x[93] = 4'd5; grid_y[93] = 4'd4;
        grid_x[94] = 4'd10; grid_y[94] = 4'd10;
        grid_x[95] = 4'd8; grid_y[95] = 4'd12;
        grid_x[96] = 4'd4; grid_y[96] = 4'd3;
        grid_x[97] = 4'd10; grid_y[97] = 4'd7;
        grid_x[98] = 4'd12; grid_y[98] = 4'd2;
        grid_x[99] = 4'd3; grid_y[99] = 4'd1;
        grid_x[100] = 4'd6; grid_y[100] = 4'd0;
        grid_x[101] = 4'd11; grid_y[101] = 4'd14;
        grid_x[102] = 4'd6; grid_y[102] = 4'd3;
        grid_x[103] = 4'd13; grid_y[103] = 4'd0;
        grid_x[104] = 4'd1; grid_y[104] = 4'd11;
        grid_x[105] = 4'd13; grid_y[105] = 4'd3;
        grid_x[106] = 4'd13; grid_y[106] = 4'd14;
        grid_x[107] = 4'd12; grid_y[107] = 4'd1;
        grid_x[108] = 4'd8; grid_y[108] = 4'd4;
        grid_x[109] = 4'd2; grid_y[109] = 4'd13;
        grid_x[110] = 4'd11; grid_y[110] = 4'd4;
        grid_x[111] = 4'd4; grid_y[111] = 4'd11;
        grid_x[112] = 4'd14; grid_y[112] = 4'd8;
        grid_x[113] = 4'd1; grid_y[113] = 4'd5;
        grid_x[114] = 4'd10; grid_y[114] = 4'd0;
        grid_x[115] = 4'd6; grid_y[115] = 4'd12;
        grid_x[116] = 4'd0; grid_y[116] = 4'd11;
        grid_x[117] = 4'd5; grid_y[117] = 4'd5;
        grid_x[118] = 4'd0; grid_y[118] = 4'd13;
        grid_x[119] = 4'd12; grid_y[119] = 4'd13;
        grid_x[120] = 4'd5; grid_y[120] = 4'd3;
        grid_x[121] = 4'd6; grid_y[121] = 4'd11;
        grid_x[122] = 4'd3; grid_y[122] = 4'd4;
        grid_x[123] = 4'd5; grid_y[123] = 4'd8;
        grid_x[124] = 4'd6; grid_y[124] = 4'd1;
        grid_x[125] = 4'd12; grid_y[125] = 4'd12;
        grid_x[126] = 4'd12; grid_y[126] = 4'd14;
        grid_x[127] = 4'd3; grid_y[127] = 4'd14;
        grid_x[128] = 4'd2; grid_y[128] = 4'd2;
        grid_x[129] = 4'd2; grid_y[129] = 4'd0;
        grid_x[130] = 4'd3; grid_y[130] = 4'd6;
        grid_x[131] = 4'd0; grid_y[131] = 4'd9;
        grid_x[132] = 4'd1; grid_y[132] = 4'd12;
        grid_x[133] = 4'd7; grid_y[133] = 4'd1;
        grid_x[134] = 4'd1; grid_y[134] = 4'd9;
        grid_x[135] = 4'd4; grid_y[135] = 4'd7;
        grid_x[136] = 4'd7; grid_y[136] = 4'd11;
        grid_x[137] = 4'd13; grid_y[137] = 4'd9;
        grid_x[138] = 4'd0; grid_y[138] = 4'd14;
        grid_x[139] = 4'd9; grid_y[139] = 4'd6;
        grid_x[140] = 4'd10; grid_y[140] = 4'd9;
        grid_x[141] = 4'd1; grid_y[141] = 4'd0;
        grid_x[142] = 4'd14; grid_y[142] = 4'd14;
        grid_x[143] = 4'd0; grid_y[143] = 4'd8;
        grid_x[144] = 4'd8; grid_y[144] = 4'd7;
        grid_x[145] = 4'd3; grid_y[145] = 4'd7;
        grid_x[146] = 4'd3; grid_y[146] = 4'd10;
        grid_x[147] = 4'd9; grid_y[147] = 4'd1;
        grid_x[148] = 4'd0; grid_y[148] = 4'd0;
        grid_x[149] = 4'd7; grid_y[149] = 4'd0;
        grid_x[150] = 4'd11; grid_y[150] = 4'd13;
        grid_x[151] = 4'd10; grid_y[151] = 4'd6;
        grid_x[152] = 4'd3; grid_y[152] = 4'd0;
        grid_x[153] = 4'd10; grid_y[153] = 4'd1;
        grid_x[154] = 4'd4; grid_y[154] = 4'd10;
        grid_x[155] = 4'd1; grid_y[155] = 4'd4;
        grid_x[156] = 4'd6; grid_y[156] = 4'd10;
        grid_x[157] = 4'd13; grid_y[157] = 4'd12;
        grid_x[158] = 4'd3; grid_y[158] = 4'd9;
        grid_x[159] = 4'd0; grid_y[159] = 4'd6;
        grid_x[160] = 4'd12; grid_y[160] = 4'd9;
        grid_x[161] = 4'd11; grid_y[161] = 4'd5;
        grid_x[162] = 4'd14; grid_y[162] = 4'd9;
        grid_x[163] = 4'd5; grid_y[163] = 4'd1;
        grid_x[164] = 4'd10; grid_y[164] = 4'd12;
        grid_x[165] = 4'd12; grid_y[165] = 4'd5;
        grid_x[166] = 4'd4; grid_y[166] = 4'd2;
        grid_x[167] = 4'd1; grid_y[167] = 4'd10;
        grid_x[168] = 4'd14; grid_y[168] = 4'd5;
        grid_x[169] = 4'd2; grid_y[169] = 4'd9;
        grid_x[170] = 4'd4; grid_y[170] = 4'd5;
        grid_x[171] = 4'd9; grid_y[171] = 4'd10;
        grid_x[172] = 4'd1; grid_y[172] = 4'd2;
        grid_x[173] = 4'd8; grid_y[173] = 4'd2;
        grid_x[174] = 4'd2; grid_y[174] = 4'd12;
        grid_x[175] = 4'd14; grid_y[175] = 4'd6;
        grid_x[176] = 4'd7; grid_y[176] = 4'd6;
        grid_x[177] = 4'd2; grid_y[177] = 4'd7;
        grid_x[178] = 4'd5; grid_y[178] = 4'd13;
        grid_x[179] = 4'd13; grid_y[179] = 4'd11;
        grid_x[180] = 4'd7; grid_y[180] = 4'd3;
        grid_x[181] = 4'd10; grid_y[181] = 4'd8;
        grid_x[182] = 4'd3; grid_y[182] = 4'd8;
        grid_x[183] = 4'd9; grid_y[183] = 4'd3;
        grid_x[184] = 4'd6; grid_y[184] = 4'd2;
        grid_x[185] = 4'd1; grid_y[185] = 4'd6;
        grid_x[186] = 4'd9; grid_y[186] = 4'd13;
        grid_x[187] = 4'd0; grid_y[187] = 4'd1;
        grid_x[188] = 4'd14; grid_y[188] = 4'd7;
        grid_x[189] = 4'd12; grid_y[189] = 4'd6;
        grid_x[190] = 4'd7; grid_y[190] = 4'd14;
        grid_x[191] = 4'd11; grid_y[191] = 4'd9;
        grid_x[192] = 4'd7; grid_y[192] = 4'd2;
        grid_x[193] = 4'd6; grid_y[193] = 4'd6;
        grid_x[194] = 4'd4; grid_y[194] = 4'd12;
        grid_x[195] = 4'd10; grid_y[195] = 4'd14;
        grid_x[196] = 4'd10; grid_y[196] = 4'd13;
        grid_x[197] = 4'd7; grid_y[197] = 4'd12;
        grid_x[198] = 4'd0; grid_y[198] = 4'd2;
        grid_x[199] = 4'd14; grid_y[199] = 4'd0;
        grid_x[200] = 4'd9; grid_y[200] = 4'd2;
        grid_x[201] = 4'd5; grid_y[201] = 4'd2;
        grid_x[202] = 4'd0; grid_y[202] = 4'd7;
        grid_x[203] = 4'd2; grid_y[203] = 4'd3;
        grid_x[204] = 4'd1; grid_y[204] = 4'd8;
        grid_x[205] = 4'd13; grid_y[205] = 4'd1;
        grid_x[206] = 4'd5; grid_y[206] = 4'd0;
        grid_x[207] = 4'd1; grid_y[207] = 4'd14;
        grid_x[208] = 4'd6; grid_y[208] = 4'd4;
        grid_x[209] = 4'd6; grid_y[209] = 4'd13;
        grid_x[210] = 4'd7; grid_y[210] = 4'd9;
        grid_x[211] = 4'd5; grid_y[211] = 4'd10;
        grid_x[212] = 4'd8; grid_y[212] = 4'd11;
        grid_x[213] = 4'd12; grid_y[213] = 4'd0;
        grid_x[214] = 4'd0; grid_y[214] = 4'd10;
        grid_x[215] = 4'd2; grid_y[215] = 4'd14;
        grid_x[216] = 4'd10; grid_y[216] = 4'd3;
        grid_x[217] = 4'd4; grid_y[217] = 4'd4;
        grid_x[218] = 4'd1; grid_y[218] = 4'd3;
        grid_x[219] = 4'd9; grid_y[219] = 4'd8;
        grid_x[220] = 4'd5; grid_y[220] = 4'd7;
        grid_x[221] = 4'd5; grid_y[221] = 4'd12;
        grid_x[222] = 4'd0; grid_y[222] = 4'd4;
        grid_x[223] = 4'd14; grid_y[223] = 4'd13;
        grid_x[224] = 4'd10; grid_y[224] = 4'd5; 

        //first spawn position.
        spawnPositionX = grid_x[0];
        spawnPositionY = grid_y[0];
    end

    always @(posedge CLOCK_50) begin
        
        if (xySelector > 223) begin
            //using blocking assignment
            xySelector <= 0;
        end  

        if ((spawnPositionX == snakePositionX) && (spawnPositionY == snakePositionY)) begin
            
            snakeLength <= snakeLength + 1;
            spawnPositionX <= grid_x[xySelector];
            spawnPositionY <= grid_y[xySelector];

            //
            //takes the last two bits of xySelector, if its 10 its fast the game, 11 is slow
            if (xySelector[1:0] == 2'b10) begin
                gameClockSelect <= 2;
            end
            else if (xySelector[1:0] == 2'b11) begin
                gameClockSelect <=1;
            end            
            else gameClockSelect <=0;
            
				//incrementing
            xySelector <= xySelector + 1;
            
				//COLOUR
            //takes the last two bits of xySelector, if its 10 its fast the game, 11 is slow
            if (xySelector[1:0] == 2'b01) begin
                itemColour <= 3'b101;
            end
            else if (xySelector[1:0] == 2'b10) begin
                itemColour <= 3'b100;
            end
            else itemColour <= 3'b010;
            
            
        end
    end 

endmodule
